library ieee;
use ieee.std_logic_1164.all;

entity HamsterBall is
port(
	clk_0,reset,datain,clkin: in std_logic;
	hs,vs: out STD_LOGIC; 
	r,g,b: out STD_LOGIC_vector(2 downto 0)
);
end HamsterBall;

architecture arc of HamsterBall is

component vga640480 is
	 port(
			address		:	  out STD_LOGIC_VECTOR(15 DOWNTO 0);
			reset       :     in  STD_LOGIC;
			clk50       :	  out std_logic; 
			qRGB		:	  in STD_LOGIC_VECTOR(8 downto 0);
			clk_0       :     in  STD_LOGIC; --50Mʱ������
			hs,vs       :     out STD_LOGIC; --��ͬ������ͬ���ź�
			r,g,b       :     out STD_LOGIC_vector(2 downto 0);
			wkey		:     in STD_LOGIC
	  );
end component;

COMPONENT mymap IS
	PORT
	(
		address		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		clock		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (8 DOWNTO 0)
	);
END COMPONENT mymap;

component top is
port(
	datain,clkin,fclk,rst_in: in std_logic;
	wkey:out std_logic
);
END component;

signal address_tmp: std_logic_vector(15 downto 0);
signal clk50: std_logic;
--signal q_red, q_green, q_blue: std_logic_vector(2 downto 0);
signal q_rgb: std_logic_vector(8 downto 0);
signal wkey: std_logic;


begin

u1: vga640480 port map(
						address=>address_tmp, 
						reset=>reset, 
						clk50=>clk50, 
						qRGB=>q_rgb,
						clk_0=>clk_0, 
						hs=>hs, vs=>vs, 
						r=>r, g=>g, b=>b,
						wkey => wkey
					);
--u2: red port map(	
--						address=>address_tmp, 
--						clock=>clk50, 
--						q=>q_red
--					);
--u3: green port map(	
--						address=>address_tmp, 
--						clock=>clk50, 
--						q=>q_green
--					);
--u4: blue port map(	
--						address=>address_tmp, 
--						clock=>clk50, 
--						q=>q_blue
--					);
u6: mymap port map(
						address=>address_tmp, 
						clock=>clk50, 
						q=>q_rgb
				  );
u5: top port map(datain,clkin,clk_0,reset,wkey);
end arc;